// setup test file
